  localparam [31:0] ADD                = 32'b0000000??????????000?????0110011;
  localparam [31:0] ADDI               = 32'b?????????????????000?????0010011;
  localparam [31:0] AND                = 32'b0000000??????????111?????0110011;
  localparam [31:0] ANDI               = 32'b?????????????????111?????0010011;
  localparam [31:0] AUIPC              = 32'b?????????????????????????0010111;
  localparam [31:0] BEQ                = 32'b?????????????????000?????1100011;
  localparam [31:0] BGE                = 32'b?????????????????101?????1100011;
  localparam [31:0] BGEU               = 32'b?????????????????111?????1100011;
  localparam [31:0] BLT                = 32'b?????????????????100?????1100011;
  localparam [31:0] BLTU               = 32'b?????????????????110?????1100011;
  localparam [31:0] BNE                = 32'b?????????????????001?????1100011;
  localparam [31:0] EBREAK             = 32'b00000000000100000000000001110011;
  localparam [31:0] ECALL              = 32'b00000000000000000000000001110011;
  localparam [31:0] FENCE              = 32'b?????????????????000?????0001111;
  localparam [31:0] JAL                = 32'b?????????????????????????1101111;
  localparam [31:0] JALR               = 32'b?????????????????000?????1100111;
  localparam [31:0] LB                 = 32'b?????????????????000?????0000011;
  localparam [31:0] LBU                = 32'b?????????????????100?????0000011;
  localparam [31:0] LH                 = 32'b?????????????????001?????0000011;
  localparam [31:0] LHU                = 32'b?????????????????101?????0000011;
  localparam [31:0] LUI                = 32'b?????????????????????????0110111;
  localparam [31:0] LW                 = 32'b?????????????????010?????0000011;
  localparam [31:0] OR                 = 32'b0000000??????????110?????0110011;
  localparam [31:0] ORI                = 32'b?????????????????110?????0010011;
  localparam [31:0] SB                 = 32'b?????????????????000?????0100011;
  localparam [31:0] SH                 = 32'b?????????????????001?????0100011;
  localparam [31:0] SLL                = 32'b0000000??????????001?????0110011;
  localparam [31:0] SLLI               = 32'b0000000??????????001?????0010011;
  localparam [31:0] SLT                = 32'b0000000??????????010?????0110011;
  localparam [31:0] SLTI               = 32'b?????????????????010?????0010011;
  localparam [31:0] SLTIU              = 32'b?????????????????011?????0010011;
  localparam [31:0] SLTU               = 32'b0000000??????????011?????0110011;
  localparam [31:0] SRA                = 32'b0100000??????????101?????0110011;
  localparam [31:0] SRAI               = 32'b0100000??????????101?????0010011;
  localparam [31:0] SRL                = 32'b0000000??????????101?????0110011;
  localparam [31:0] SRLI               = 32'b0000000??????????101?????0010011;
  localparam [31:0] SUB                = 32'b0100000??????????000?????0110011;
  localparam [31:0] SW                 = 32'b?????????????????010?????0100011;
  localparam [31:0] XOR                = 32'b0000000??????????100?????0110011;
  localparam [31:0] XORI               = 32'b?????????????????100?????0010011;
